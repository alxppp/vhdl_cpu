package cpu_subprogram_pack_alex is

use WORK.cpu_defs_pack.all;
use WORK.bit_vector_natural_pack.all;

end cpu_subprogram_pack_alex;

package body cpu_subprogram_pack_alex is

end cpu_subprogram_pack_alex;
