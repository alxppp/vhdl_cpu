package cpu_subprogram_pack_robert is

use WORK.cpu_defs_pack.all;
use WORK.bit_vector_natural_pack.all;

end cpu_subprogram_pack_robert;

package body cpu_subprogram_pack_robert is


end cpu_subprogram_pack_robert;