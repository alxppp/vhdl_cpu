package cpu_subprogram_pack_max is





end cpu_subprogram_pack_max;


package body cpu_subprogram_pack_max is




end cpu_subprogram_pack_max;